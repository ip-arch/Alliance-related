* Spice description of pvssck2_sp
* Spice driver version 4802095
* Date ( dd/mm/yyyy hh:mm:ss ): 11/12/2016 at 17:45:24

* INTERF ck cko vdd vss 


.subckt pvssck2_sp 4 3 5 6 
* NET 3 = cko
* NET 4 = ck
* NET 5 = vdd
* NET 6 = vss
Mtr_00019 3 2 5 5 tp L=2U W=61.5U AS=430.5P AD=430.5P PS=137U PD=137U 
Mtr_00018 5 2 3 5 tp L=2U W=61.5U AS=430.5P AD=430.5P PS=137U PD=137U 
Mtr_00017 3 2 5 5 tp L=2U W=61.5U AS=430.5P AD=430.5P PS=137U PD=137U 
Mtr_00016 5 2 3 5 tp L=2U W=61.5U AS=430.5P AD=430.5P PS=137U PD=137U 
Mtr_00015 3 2 5 5 tp L=2U W=61.5U AS=430.5P AD=430.5P PS=137U PD=137U 
Mtr_00014 5 2 3 5 tp L=2U W=61.5U AS=430.5P AD=430.5P PS=137U PD=137U 
Mtr_00013 5 2 3 5 tp L=2U W=61.5U AS=430.5P AD=430.5P PS=137U PD=137U 
Mtr_00012 5 2 3 5 tp L=2U W=61.5U AS=430.5P AD=430.5P PS=137U PD=137U 
Mtr_00011 5 4 2 5 tp L=2U W=49U AS=343P AD=343P PS=112U PD=112U 
Mtr_00010 5 2 3 5 tp L=2U W=49U AS=343P AD=343P PS=112U PD=112U 
Mtr_00009 3 2 5 5 tp L=2U W=49U AS=343P AD=343P PS=112U PD=112U 
Mtr_00008 5 2 3 5 tp L=2U W=49U AS=343P AD=343P PS=112U PD=112U 
Mtr_00007 3 2 5 5 tp L=2U W=49U AS=343P AD=343P PS=112U PD=112U 
Mtr_00006 5 4 2 5 tp L=2U W=136.5U AS=955.5P AD=955.5P PS=287U PD=287U 
Mtr_00005 3 2 6 6 tn L=2U W=61.5U AS=430.5P AD=430.5P PS=137U PD=137U 
Mtr_00004 6 2 3 6 tn L=2U W=61.5U AS=430.5P AD=430.5P PS=137U PD=137U 
Mtr_00003 3 2 6 6 tn L=2U W=61.5U AS=430.5P AD=430.5P PS=137U PD=137U 
Mtr_00002 6 2 3 6 tn L=2U W=61.5U AS=430.5P AD=430.5P PS=137U PD=137U 
Mtr_00001 6 4 2 6 tn L=2U W=61.5U AS=430.5P AD=430.5P PS=137U PD=137U 
.ends pvssck2_sp

